* WARNING : please consider following remarks before usage
*
* 1) All models are a tradeoff between accuracy and complexity (ie. simulation 
*    time).
* 2) Macromodels are not a substitute to breadboarding, they rather confirm the
*    validity of a design approach and help to select surrounding component values.
*
* 3) A macromodel emulates the NOMINAL performance of a TYPICAL device within 
*    SPECIFIED OPERATING CONDITIONS (ie. temperature, supply voltage, etc.).
*    Thus the macromodel is often not as exhaustive as the datasheet, its goal
*    is to illustrate the main parameters of the product.
*
* 4) Data issued from macromodels used outside of its specified conditions
*    (Vcc, Temperature, etc) or even worse: outside of the device operating 
*    conditions (Vcc, Vicm, etc) are not reliable in any way.


** Macanal, Analog macromodels generator, v.1.0
** J. REMY, SGS THOMSON, ANACA Grenoble, Aug. 1992.
** Standard Linear Ics Macromodels, 1993. 
** CONNECTIONS :
* 1 INVERTING INPUT
* 2 NON-INVERTING INPUT
* 3 OUTPUT
* 4 POSITIVE POWER SUPPLY
* 5 NEGATIVE POWER SUPPLY
.SUBCKT LM101 1 3 2 4 5 (analog)
********************************************************
.MODEL MDTH D IS=1E-8 KF=1.025862E-15 CJO=10F
* INPUT STAGE
CIP 2 5 1.000000E-12
CIN 1 5 1.000000E-12
EIP 10 5 2 5 1
EIN 16 5 1 5 1
RIP 10 11 1.625000E+01
RIN 15 16 1.625000E+01
RIS 11 15 7.476714E+01
DIP 11 12 MDTH 400E-12
DIN 15 14 MDTH 400E-12
VOFP 12 13 DC 0.000000E+00
VOFN 13 14 DC 0
IPOL 13 5 1.600000E-05
CPS 11 15 2.5E-09
DINN 17 13 MDTH 400E-12
VIN 17 5 0.000000e+00
DINR 15 18 MDTH 400E-12
VIP 4 18 0.000000E+00
FCP 4 5 VOFP 1.115000E+02
FCN 5 4 VOFN 1.115000E+02
FIBP 2 5 VOFP 1.875000E-04
FIBN 5 1 VOFN 1.875000E-04
* AMPLIFYING STAGE
FIP 5 19 VOFP 9.375000E+02
FIN 5 19 VOFN 9.375000E+02
RG1 19 5 9.981802E+05
RG2 19 4 9.981802E+05
CC 19 29 3.000000E-08
HZTP 30 29 VOFP 5.535733E+02
HZTN  5 30 VOFN 5.535733E+02
DOPM 19 22 MDTH 400E-12
DONM 21 19 MDTH 400E-12
HOPM 22 28 VOUT 5.000000E+03
VIPM 28 4 1.500000E+02
HONM 21 27 VOUT 5.000000E+03
VINM 5 27 1.500000E+02
EOUT 26 23 19 5 1
VOUT 23 5 0
ROUT 26 3 200
COUT 3 5 1.000000E-12
DOP 19 25 MDTH 400E-12
VOP 4 25 1.480450E+00
DON 24 19 MDTH 400E-12
VON 24 5 1.480450E+00
.ENDS